module tb();
reg signed [31:0] L1;
reg signed [31:0] L2;
reg signed [31:0] L3;
reg signed [31:0] L4;
reg signed [31:0] L5;
reg signed [31:0] L6;
reg signed [31:0] L7;
reg signed [31:0] L8;
reg signed [31:0] L9;
reg signed [31:0] L10;
reg signed [31:0] L11;
reg signed [31:0] L12;
reg signed [31:0] L13;
reg signed [31:0] L14;
reg signed [31:0] L15;
reg signed [31:0] L16;
reg signed [31:0] L17;
reg signed [31:0] L18;
reg signed [31:0] L19;
reg signed [31:0] L20;
reg signed [31:0] L21;
reg signed [31:0] L22;
reg signed [31:0] L23;
reg signed [31:0] L24;
reg signed [31:0] L25;
reg signed [31:0] L26;
reg signed [31:0] L27;
reg signed [31:0] L28;
reg signed [31:0] L29;
reg signed [31:0] L30;
reg signed [31:0] L31;
reg signed [31:0] L32;
reg signed [31:0] L33;
reg signed [31:0] L34;
reg signed [31:0] L35;
reg signed [31:0] L36;
reg signed [31:0] L37;
reg signed [31:0] L38;
reg signed [31:0] L39;
reg signed [31:0] L40;
reg signed [31:0] L41;
reg signed [31:0] L42;
reg signed [31:0] L43;
reg signed [31:0] L44;
reg signed [31:0] L45;
reg signed [31:0] L46;
reg signed [31:0] L47;
reg signed [31:0] L48;
reg signed [31:0] L49;
reg signed [31:0] L50;
reg signed [31:0] L51;
reg signed [31:0] L52;
reg signed [31:0] L53;
reg signed [31:0] L54;
reg signed [31:0] L55;
reg signed [31:0] L56;
reg signed [31:0] L57;
reg signed [31:0] L58;
reg signed [31:0] L59;
reg signed [31:0] L60;
reg signed [31:0] L61;
reg signed [31:0] L62;
reg signed [31:0] L63;
reg signed [31:0] L64;
reg signed [31:0] L65;
reg signed [31:0] L66;
reg signed [31:0] L67;
reg signed [31:0] L68;
reg signed [31:0] L69;
reg signed [31:0] L70;
reg signed [31:0] L71;
reg signed [31:0] L72;
reg signed [31:0] L73;
reg signed [31:0] L74;
reg signed [31:0] L75;
reg signed [31:0] L76;
reg signed [31:0] L77;
reg signed [31:0] L78;
reg signed [31:0] L79;
reg signed [31:0] L80;
reg signed [31:0] L81;
reg signed [31:0] L82;
reg signed [31:0] L83;
reg signed [31:0] L84;
reg signed [31:0] L85;
reg signed [31:0] L86;
reg signed [31:0] L87;
reg signed [31:0] L88;
reg signed [31:0] L89;
reg signed [31:0] L90;
reg signed [31:0] L91;
reg signed [31:0] L92;
reg signed [31:0] L93;
reg signed [31:0] L94;
reg signed [31:0] L95;
reg signed [31:0] L96;
reg signed [31:0] L97;
reg signed [31:0] L98;
reg signed [31:0] L99;
reg signed [31:0] L100;
reg signed [31:0] L101;
reg signed [31:0] L102;
reg signed [31:0] L103;
reg signed [31:0] L104;
reg signed [31:0] L105;
reg signed [31:0] L106;
reg signed [31:0] L107;
reg signed [31:0] L108;
reg signed [31:0] L109;
reg signed [31:0] L110;
reg signed [31:0] L111;
reg signed [31:0] L112;
reg signed [31:0] L113;
reg signed [31:0] L114;
reg signed [31:0] L115;
reg signed [31:0] L116;
reg signed [31:0] L117;
reg signed [31:0] L118;
reg signed [31:0] L119;
reg signed [31:0] L120;
reg signed [31:0] L121;
reg signed [31:0] L122;
reg signed [31:0] L123;
reg signed [31:0] L124;
reg signed [31:0] L125;
reg signed [31:0] L126;
reg signed [31:0] L127;
reg signed [31:0] L128;
reg signed [31:0] L129;
reg signed [31:0] L130;
reg signed [31:0] L131;
reg signed [31:0] L132;
reg signed [31:0] L133;
reg signed [31:0] L134;
reg signed [31:0] L135;
reg signed [31:0] L136;
reg signed [31:0] L137;
reg signed [31:0] L138;
reg signed [31:0] L139;
reg signed [31:0] L140;
reg signed [31:0] L141;
reg signed [31:0] L142;
reg signed [31:0] L143;
reg signed [31:0] L144;
reg signed [31:0] L145;
reg signed [31:0] L146;
reg signed [31:0] L147;
reg signed [31:0] L148;
reg signed [31:0] L149;
reg signed [31:0] L150;
reg signed [31:0] L151;
reg signed [31:0] L152;
reg signed [31:0] L153;
reg signed [31:0] L154;
reg signed [31:0] L155;
reg signed [31:0] L156;
reg signed [31:0] L157;
reg signed [31:0] L158;
reg signed [31:0] L159;
reg signed [31:0] L160;
reg signed [31:0] L161;
reg signed [31:0] L162;
reg signed [31:0] L163;
reg signed [31:0] L164;
reg signed [31:0] L165;
reg signed [31:0] L166;
reg signed [31:0] L167;
reg signed [31:0] L168;
reg signed [31:0] L169;
reg signed [31:0] L170;
reg signed [31:0] L171;
reg signed [31:0] L172;
reg signed [31:0] L173;
reg signed [31:0] L174;
reg signed [31:0] L175;
reg signed [31:0] L176;
reg signed [31:0] L177;
reg signed [31:0] L178;
reg signed [31:0] L179;
reg signed [31:0] L180;
reg signed [31:0] L181;
reg signed [31:0] L182;
reg signed [31:0] L183;
reg signed [31:0] L184;
reg signed [31:0] L185;
reg signed [31:0] L186;
reg signed [31:0] L187;
reg signed [31:0] L188;
reg signed [31:0] L189;
reg signed [31:0] L190;
reg signed [31:0] L191;
reg signed [31:0] L192;
reg signed [31:0] L193;
reg signed [31:0] L194;
reg signed [31:0] L195;
reg signed [31:0] L196;
reg signed [31:0] L197;
reg signed [31:0] L198;
reg signed [31:0] L199;
reg signed [31:0] L200;
reg signed [31:0] L201;
reg signed [31:0] L202;
reg signed [31:0] L203;
reg signed [31:0] L204;
reg signed [31:0] L205;
reg signed [31:0] L206;
reg signed [31:0] L207;
reg signed [31:0] L208;
reg signed [31:0] L209;
reg signed [31:0] L210;
reg signed [31:0] L211;
reg signed [31:0] L212;
reg signed [31:0] L213;
reg signed [31:0] L214;
reg signed [31:0] L215;
reg signed [31:0] L216;
reg signed [31:0] L217;
reg signed [31:0] L218;
reg signed [31:0] L219;
reg signed [31:0] L220;
reg signed [31:0] L221;
reg signed [31:0] L222;
reg signed [31:0] L223;
reg signed [31:0] L224;
reg signed [31:0] L225;
reg signed [31:0] L226;
reg signed [31:0] L227;
reg signed [31:0] L228;
reg signed [31:0] L229;
reg signed [31:0] L230;
reg signed [31:0] L231;
reg signed [31:0] L232;
reg signed [31:0] L233;
reg signed [31:0] L234;
reg signed [31:0] L235;
reg signed [31:0] L236;
reg signed [31:0] L237;
reg signed [31:0] L238;
reg signed [31:0] L239;
reg signed [31:0] L240;
reg signed [31:0] L241;
reg signed [31:0] L242;
reg signed [31:0] L243;
reg signed [31:0] L244;
reg signed [31:0] L245;
reg signed [31:0] L246;
reg signed [31:0] L247;
reg signed [31:0] L248;
reg signed [31:0] L249;
reg signed [31:0] L250;
reg signed [31:0] L251;
reg signed [31:0] L252;
reg signed [31:0] L253;
reg signed [31:0] L254;
reg signed [31:0] L255;
reg signed [31:0] L256;
reg signed [31:0] L257;
reg signed [31:0] L258;
reg signed [31:0] L259;
reg signed [31:0] L260;
reg signed [31:0] L261;
reg signed [31:0] L262;
reg signed [31:0] L263;
reg signed [31:0] L264;
reg signed [31:0] L265;
reg signed [31:0] L266;
reg signed [31:0] L267;
reg signed [31:0] L268;
reg signed [31:0] L269;
reg signed [31:0] L270;
reg signed [31:0] L271;
reg signed [31:0] L272;
reg signed [31:0] L273;
reg signed [31:0] L274;
reg signed [31:0] L275;
reg signed [31:0] L276;
reg signed [31:0] L277;
reg signed [31:0] L278;
reg signed [31:0] L279;
reg signed [31:0] L280;
reg signed [31:0] L281;
reg signed [31:0] L282;
reg signed [31:0] L283;
reg signed [31:0] L284;
reg signed [31:0] L285;
reg signed [31:0] L286;
reg signed [31:0] L287;
reg signed [31:0] L288;
reg signed [31:0] L289;
reg signed [31:0] L290;
reg signed [31:0] L291;
reg signed [31:0] L292;
reg signed [31:0] L293;
reg signed [31:0] L294;
reg signed [31:0] L295;
reg signed [31:0] L296;
reg signed [31:0] L297;
reg signed [31:0] L298;
reg signed [31:0] L299;
reg signed [31:0] L300;
reg signed [31:0] L301;
reg signed [31:0] L302;
reg signed [31:0] L303;
reg signed [31:0] L304;
reg signed [31:0] L305;
reg signed [31:0] L306;
reg signed [31:0] L307;
reg signed [31:0] L308;
reg signed [31:0] L309;
reg signed [31:0] L310;
reg signed [31:0] L311;
reg signed [31:0] L312;
reg signed [31:0] L313;
reg signed [31:0] L314;
reg signed [31:0] L315;
reg signed [31:0] L316;
reg signed [31:0] L317;
reg signed [31:0] L318;
reg signed [31:0] L319;
reg signed [31:0] L320;
reg signed [31:0] L321;
reg signed [31:0] L322;
reg signed [31:0] L323;
reg signed [31:0] L324;
reg signed [31:0] L325;
reg signed [31:0] L326;
reg signed [31:0] L327;
reg signed [31:0] L328;
reg signed [31:0] L329;
reg signed [31:0] L330;
reg signed [31:0] L331;
reg signed [31:0] L332;
reg signed [31:0] L333;
reg signed [31:0] L334;
reg signed [31:0] L335;
reg signed [31:0] L336;
reg signed [31:0] L337;
reg signed [31:0] L338;
reg signed [31:0] L339;
reg signed [31:0] L340;
reg signed [31:0] L341;
reg signed [31:0] L342;
reg signed [31:0] L343;
reg signed [31:0] L344;
reg signed [31:0] L345;
reg signed [31:0] L346;
reg signed [31:0] L347;
reg signed [31:0] L348;
reg signed [31:0] L349;
reg signed [31:0] L350;
reg signed [31:0] L351;
reg signed [31:0] L352;
reg signed [31:0] L353;
reg signed [31:0] L354;
reg signed [31:0] L355;
reg signed [31:0] L356;
reg signed [31:0] L357;
reg signed [31:0] L358;
reg signed [31:0] L359;
reg signed [31:0] L360;
reg signed [31:0] L361;
reg signed [31:0] L362;
reg signed [31:0] L363;
reg signed [31:0] L364;
reg signed [31:0] L365;
reg signed [31:0] L366;
reg signed [31:0] L367;
reg signed [31:0] L368;
reg signed [31:0] L369;
reg signed [31:0] L370;
reg signed [31:0] L371;
reg signed [31:0] L372;
reg signed [31:0] L373;
reg signed [31:0] L374;
reg signed [31:0] L375;
reg signed [31:0] L376;
reg signed [31:0] L377;
reg signed [31:0] L378;
reg signed [31:0] L379;
reg signed [31:0] L380;
reg signed [31:0] L381;
reg signed [31:0] L382;
reg signed [31:0] L383;
reg signed [31:0] L384;
reg signed [31:0] L385;
reg signed [31:0] L386;
reg signed [31:0] L387;
reg signed [31:0] L388;
reg signed [31:0] L389;
reg signed [31:0] L390;
reg signed [31:0] L391;
reg signed [31:0] L392;
reg signed [31:0] L393;
reg signed [31:0] L394;
reg signed [31:0] L395;
reg signed [31:0] L396;
reg signed [31:0] L397;
reg signed [31:0] L398;
reg signed [31:0] L399;
reg signed [31:0] L400;
reg signed [31:0] L401;
reg signed [31:0] L402;
reg signed [31:0] L403;
reg signed [31:0] L404;
reg signed [31:0] L405;
reg signed [31:0] L406;
reg signed [31:0] L407;
reg signed [31:0] L408;
reg signed [31:0] L409;
reg signed [31:0] L410;
reg signed [31:0] L411;
reg signed [31:0] L412;
reg signed [31:0] L413;
reg signed [31:0] L414;
reg signed [31:0] L415;
reg signed [31:0] L416;
reg signed [31:0] L417;
reg signed [31:0] L418;
reg signed [31:0] L419;
reg signed [31:0] L420;
reg signed [31:0] L421;
reg signed [31:0] L422;
reg signed [31:0] L423;
reg signed [31:0] L424;
reg signed [31:0] L425;
reg signed [31:0] L426;
reg signed [31:0] L427;
reg signed [31:0] L428;
reg signed [31:0] L429;
reg signed [31:0] L430;
reg signed [31:0] L431;
reg signed [31:0] L432;
reg signed [31:0] L433;
reg signed [31:0] L434;
reg signed [31:0] L435;
reg signed [31:0] L436;
reg signed [31:0] L437;
reg signed [31:0] L438;
reg signed [31:0] L439;
reg signed [31:0] L440;
reg signed [31:0] L441;
reg signed [31:0] L442;
reg signed [31:0] L443;
reg signed [31:0] L444;
reg signed [31:0] L445;
reg signed [31:0] L446;
reg signed [31:0] L447;
reg signed [31:0] L448;
reg signed [31:0] L449;
reg signed [31:0] L450;
reg signed [31:0] L451;
reg signed [31:0] L452;
reg signed [31:0] L453;
reg signed [31:0] L454;
reg signed [31:0] L455;
reg signed [31:0] L456;
reg signed [31:0] L457;
reg signed [31:0] L458;
reg signed [31:0] L459;
reg signed [31:0] L460;
reg signed [31:0] L461;
reg signed [31:0] L462;
reg signed [31:0] L463;
reg signed [31:0] L464;
reg signed [31:0] L465;
reg signed [31:0] L466;
reg signed [31:0] L467;
reg signed [31:0] L468;
reg signed [31:0] L469;
reg signed [31:0] L470;
reg signed [31:0] L471;
reg signed [31:0] L472;
reg signed [31:0] L473;
reg signed [31:0] L474;
reg signed [31:0] L475;
reg signed [31:0] L476;
reg signed [31:0] L477;
reg signed [31:0] L478;
reg signed [31:0] L479;
reg signed [31:0] L480;
reg signed [31:0] L481;
reg signed [31:0] L482;
reg signed [31:0] L483;
reg signed [31:0] L484;
reg signed [31:0] L485;
reg signed [31:0] L486;
reg signed [31:0] L487;
reg signed [31:0] L488;
reg signed [31:0] L489;
reg signed [31:0] L490;
reg signed [31:0] L491;
reg signed [31:0] L492;
reg signed [31:0] L493;
reg signed [31:0] L494;
reg signed [31:0] L495;
reg signed [31:0] L496;
reg signed [31:0] L497;
reg signed [31:0] L498;
reg signed [31:0] L499;
reg signed [31:0] L500;
reg signed [31:0] L501;
reg signed [31:0] L502;
reg signed [31:0] L503;
reg signed [31:0] L504;
reg signed [31:0] L505;
reg signed [31:0] L506;
reg signed [31:0] L507;
reg signed [31:0] L508;
reg signed [31:0] L509;
reg signed [31:0] L510;
reg signed [31:0] L511;
reg signed [31:0] L512;
reg signed [31:0] L513;
reg signed [31:0] L514;
reg signed [31:0] L515;
reg signed [31:0] L516;
reg signed [31:0] L517;
reg signed [31:0] L518;
reg signed [31:0] L519;
reg signed [31:0] L520;
reg signed [31:0] L521;
reg signed [31:0] L522;
reg signed [31:0] L523;
reg signed [31:0] L524;
reg signed [31:0] L525;
reg signed [31:0] L526;
reg signed [31:0] L527;
reg signed [31:0] L528;
reg signed [31:0] L529;
reg signed [31:0] L530;
reg signed [31:0] L531;
reg signed [31:0] L532;
reg signed [31:0] L533;
reg signed [31:0] L534;
reg signed [31:0] L535;
reg signed [31:0] L536;
reg signed [31:0] L537;
reg signed [31:0] L538;
reg signed [31:0] L539;
reg signed [31:0] L540;
reg signed [31:0] L541;
reg signed [31:0] L542;
reg signed [31:0] L543;
reg signed [31:0] L544;
reg signed [31:0] L545;
reg signed [31:0] L546;
reg signed [31:0] L547;
reg signed [31:0] L548;
reg signed [31:0] L549;
reg signed [31:0] L550;
reg signed [31:0] L551;
reg signed [31:0] L552;
reg signed [31:0] L553;
reg signed [31:0] L554;
reg signed [31:0] L555;
reg signed [31:0] L556;
reg signed [31:0] L557;
reg signed [31:0] L558;
reg signed [31:0] L559;
reg signed [31:0] L560;
reg signed [31:0] L561;
reg signed [31:0] L562;
reg signed [31:0] L563;
reg signed [31:0] L564;
reg signed [31:0] L565;
reg signed [31:0] L566;
reg signed [31:0] L567;
reg signed [31:0] L568;
reg signed [31:0] L569;
reg signed [31:0] L570;
reg signed [31:0] L571;
reg signed [31:0] L572;
reg signed [31:0] L573;
reg signed [31:0] L574;
reg signed [31:0] L575;
reg signed [31:0] L576;
wire [575:0] P;
reg clk;reg rst;
LDPC_decoder_TOP LDPC1(clk,rst,L1,L2,L3,L4,L5,L6,L7,L8,L9,L10,L11,L12,L13,L14,L15,L16,L17,L18,L19,L20,L21,L22,L23,L24,L25,L26,L27,L28,L29,L30,L31,L32,L33,L34,L35,L36,L37,L38,L39,L40,L41,L42,L43,L44,L45,L46,L47,L48,L49,L50,L51,L52,L53,L54,L55,L56,L57,L58,L59,L60,L61,L62,L63,L64,L65,L66,L67,L68,L69,L70,L71,L72,L73,L74,L75,L76,L77,L78,L79,L80,L81,L82,L83,L84,L85,L86,L87,L88,L89,L90,L91,L92,L93,L94,L95,L96,L97,L98,L99,L100,L101,L102,L103,L104,L105,L106,L107,L108,L109,L110,L111,L112,L113,L114,L115,L116,L117,L118,L119,L120,L121,L122,L123,L124,L125,L126,L127,L128,L129,L130,L131,L132,L133,L134,L135,L136,L137,L138,L139,L140,L141,L142,L143,L144,L145,L146,L147,L148,L149,L150,L151,L152,L153,L154,L155,L156,L157,L158,L159,L160,L161,L162,L163,L164,L165,L166,L167,L168,L169,L170,L171,L172,L173,L174,L175,L176,L177,L178,L179,L180,L181,L182,L183,L184,L185,L186,L187,L188,L189,L190,L191,L192,L193,L194,L195,L196,L197,L198,L199,L200,L201,L202,L203,L204,L205,L206,L207,L208,L209,L210,L211,L212,L213,L214,L215,L216,L217,L218,L219,L220,L221,L222,L223,L224,L225,L226,L227,L228,L229,L230,L231,L232,L233,L234,L235,L236,L237,L238,L239,L240,L241,L242,L243,L244,L245,L246,L247,L248,L249,L250,L251,L252,L253,L254,L255,L256,L257,L258,L259,L260,L261,L262,L263,L264,L265,L266,L267,L268,L269,L270,L271,L272,L273,L274,L275,L276,L277,L278,L279,L280,L281,L282,L283,L284,L285,L286,L287,L288,L289,L290,L291,L292,L293,L294,L295,L296,L297,L298,L299,L300,L301,L302,L303,L304,L305,L306,L307,L308,L309,L310,L311,L312,L313,L314,L315,L316,L317,L318,L319,L320,L321,L322,L323,L324,L325,L326,L327,L328,L329,L330,L331,L332,L333,L334,L335,L336,L337,L338,L339,L340,L341,L342,L343,L344,L345,L346,L347,L348,L349,L350,L351,L352,L353,L354,L355,L356,L357,L358,L359,L360,L361,L362,L363,L364,L365,L366,L367,L368,L369,L370,L371,L372,L373,L374,L375,L376,L377,L378,L379,L380,L381,L382,L383,L384,L385,L386,L387,L388,L389,L390,L391,L392,L393,L394,L395,L396,L397,L398,L399,L400,L401,L402,L403,L404,L405,L406,L407,L408,L409,L410,L411,L412,L413,L414,L415,L416,L417,L418,L419,L420,L421,L422,L423,L424,L425,L426,L427,L428,L429,L430,L431,L432,L433,L434,L435,L436,L437,L438,L439,L440,L441,L442,L443,L444,L445,L446,L447,L448,L449,L450,L451,L452,L453,L454,L455,L456,L457,L458,L459,L460,L461,L462,L463,L464,L465,L466,L467,L468,L469,L470,L471,L472,L473,L474,L475,L476,L477,L478,L479,L480,L481,L482,L483,L484,L485,L486,L487,L488,L489,L490,L491,L492,L493,L494,L495,L496,L497,L498,L499,L500,L501,L502,L503,L504,L505,L506,L507,L508,L509,L510,L511,L512,L513,L514,L515,L516,L517,L518,L519,L520,L521,L522,L523,L524,L525,L526,L527,L528,L529,L530,L531,L532,L533,L534,L535,L536,L537,L538,L539,L540,L541,L542,L543,L544,L545,L546,L547,L548,L549,L550,L551,L552,L553,L554,L555,L556,L557,L558,L559,L560,L561,L562,L563,L564,L565,L566,L567,L568,L569,L570,L571,L572,L573,L574,L575,L576,P[0],P[1],P[2],P[3],P[4],P[5],P[6],P[7],P[8],P[9],P[10],P[11],P[12],P[13],P[14],P[15],P[16],P[17],P[18],P[19],P[20],P[21],P[22],P[23],P[24],P[25],P[26],P[27],P[28],P[29],P[30],P[31],P[32],P[33],P[34],P[35],P[36],P[37],P[38],P[39],P[40],P[41],P[42],P[43],P[44],P[45],P[46],P[47],P[48],P[49],P[50],P[51],P[52],P[53],P[54],P[55],P[56],P[57],P[58],P[59],P[60],P[61],P[62],P[63],P[64],P[65],P[66],P[67],P[68],P[69],P[70],P[71],P[72],P[73],P[74],P[75],P[76],P[77],P[78],P[79],P[80],P[81],P[82],P[83],P[84],P[85],P[86],P[87],P[88],P[89],P[90],P[91],P[92],P[93],P[94],P[95],P[96],P[97],P[98],P[99],P[100],P[101],P[102],P[103],P[104],P[105],P[106],P[107],P[108],P[109],P[110],P[111],P[112],P[113],P[114],P[115],P[116],P[117],P[118],P[119],P[120],P[121],P[122],P[123],P[124],P[125],P[126],P[127],P[128],P[129],P[130],P[131],P[132],P[133],P[134],P[135],P[136],P[137],P[138],P[139],P[140],P[141],P[142],P[143],P[144],P[145],P[146],P[147],P[148],P[149],P[150],P[151],P[152],P[153],P[154],P[155],P[156],P[157],P[158],P[159],P[160],P[161],P[162],P[163],P[164],P[165],P[166],P[167],P[168],P[169],P[170],P[171],P[172],P[173],P[174],P[175],P[176],P[177],P[178],P[179],P[180],P[181],P[182],P[183],P[184],P[185],P[186],P[187],P[188],P[189],P[190],P[191],P[192],P[193],P[194],P[195],P[196],P[197],P[198],P[199],P[200],P[201],P[202],P[203],P[204],P[205],P[206],P[207],P[208],P[209],P[210],P[211],P[212],P[213],P[214],P[215],P[216],P[217],P[218],P[219],P[220],P[221],P[222],P[223],P[224],P[225],P[226],P[227],P[228],P[229],P[230],P[231],P[232],P[233],P[234],P[235],P[236],P[237],P[238],P[239],P[240],P[241],P[242],P[243],P[244],P[245],P[246],P[247],P[248],P[249],P[250],P[251],P[252],P[253],P[254],P[255],P[256],P[257],P[258],P[259],P[260],P[261],P[262],P[263],P[264],P[265],P[266],P[267],P[268],P[269],P[270],P[271],P[272],P[273],P[274],P[275],P[276],P[277],P[278],P[279],P[280],P[281],P[282],P[283],P[284],P[285],P[286],P[287],P[288],P[289],P[290],P[291],P[292],P[293],P[294],P[295],P[296],P[297],P[298],P[299],P[300],P[301],P[302],P[303],P[304],P[305],P[306],P[307],P[308],P[309],P[310],P[311],P[312],P[313],P[314],P[315],P[316],P[317],P[318],P[319],P[320],P[321],P[322],P[323],P[324],P[325],P[326],P[327],P[328],P[329],P[330],P[331],P[332],P[333],P[334],P[335],P[336],P[337],P[338],P[339],P[340],P[341],P[342],P[343],P[344],P[345],P[346],P[347],P[348],P[349],P[350],P[351],P[352],P[353],P[354],P[355],P[356],P[357],P[358],P[359],P[360],P[361],P[362],P[363],P[364],P[365],P[366],P[367],P[368],P[369],P[370],P[371],P[372],P[373],P[374],P[375],P[376],P[377],P[378],P[379],P[380],P[381],P[382],P[383],P[384],P[385],P[386],P[387],P[388],P[389],P[390],P[391],P[392],P[393],P[394],P[395],P[396],P[397],P[398],P[399],P[400],P[401],P[402],P[403],P[404],P[405],P[406],P[407],P[408],P[409],P[410],P[411],P[412],P[413],P[414],P[415],P[416],P[417],P[418],P[419],P[420],P[421],P[422],P[423],P[424],P[425],P[426],P[427],P[428],P[429],P[430],P[431],P[432],P[433],P[434],P[435],P[436],P[437],P[438],P[439],P[440],P[441],P[442],P[443],P[444],P[445],P[446],P[447],P[448],P[449],P[450],P[451],P[452],P[453],P[454],P[455],P[456],P[457],P[458],P[459],P[460],P[461],P[462],P[463],P[464],P[465],P[466],P[467],P[468],P[469],P[470],P[471],P[472],P[473],P[474],P[475],P[476],P[477],P[478],P[479],P[480],P[481],P[482],P[483],P[484],P[485],P[486],P[487],P[488],P[489],P[490],P[491],P[492],P[493],P[494],P[495],P[496],P[497],P[498],P[499],P[500],P[501],P[502],P[503],P[504],P[505],P[506],P[507],P[508],P[509],P[510],P[511],P[512],P[513],P[514],P[515],P[516],P[517],P[518],P[519],P[520],P[521],P[522],P[523],P[524],P[525],P[526],P[527],P[528],P[529],P[530],P[531],P[532],P[533],P[534],P[535],P[536],P[537],P[538],P[539],P[540],P[541],P[542],P[543],P[544],P[545],P[546],P[547],P[548],P[549],P[550],P[551],P[552],P[553],P[554],P[555],P[556],P[557],P[558],P[559],P[560],P[561],P[562],P[563],P[564],P[565],P[566],P[567],P[568],P[569],P[570],P[571],P[572],P[573],P[574],P[575]);
initial begin
#0 clk =1'b0;
#0 rst = 1'b1;
#5 clk =1'b1;
#5 clk =1'b0;
#5 clk =1'b1;
#20 rst = 1'b0;
forever #5 clk = ~clk;
end
initial
begin
L1 = 32'd553;
L2 = -32'd562;
L3 = 32'd870;
L4 = 32'd398;
L5 = 32'd43;
L6 = -32'd64;
L7 = 32'd841;
L8 = 32'd609;
L9 = 32'd15;
L10 = 32'd508;
L11 = 32'd281;
L12 = 32'd524;
L13 = 32'd612;
L14 = 32'd332;
L15 = 32'd67;
L16 = 32'd1795;
L17 = -32'd282;
L18 = 32'd839;
L19 = -32'd253;
L20 = -32'd30;
L21 = 32'd952;
L22 = 32'd711;
L23 = -32'd22;
L24 = 32'd1007;
L25 = -32'd81;
L26 = 32'd622;
L27 = 32'd243;
L28 = 32'd408;
L29 = 32'd522;
L30 = 32'd1110;
L31 = 32'd428;
L32 = 32'd131;
L33 = 32'd723;
L34 = 32'd183;
L35 = -32'd609;
L36 = 32'd859;
L37 = 32'd1052;
L38 = 32'd876;
L39 = 32'd745;
L40 = 32'd379;
L41 = 32'd684;
L42 = 32'd1071;
L43 = 32'd155;
L44 = 32'd15;
L45 = 32'd785;
L46 = 32'd1119;
L47 = -32'd73;
L48 = -32'd20;
L49 = 32'd1056;
L50 = 32'd308;
L51 = 32'd821;
L52 = 32'd324;
L53 = 32'd1149;
L54 = 32'd1548;
L55 = 32'd314;
L56 = 32'd1400;
L57 = 32'd1690;
L58 = 32'd570;
L59 = -32'd173;
L60 = 32'd769;
L61 = 32'd2132;
L62 = 32'd370;
L63 = 32'd990;
L64 = 32'd911;
L65 = 32'd645;
L66 = 32'd699;
L67 = -32'd304;
L68 = 32'd1261;
L69 = 32'd243;
L70 = 32'd318;
L71 = 32'd740;
L72 = 32'd149;
L73 = 32'd344;
L74 = 32'd189;
L75 = 32'd215;
L76 = 32'd1121;
L77 = -32'd174;
L78 = -32'd558;
L79 = 32'd1163;
L80 = 32'd2030;
L81 = 32'd698;
L82 = 32'd440;
L83 = 32'd1163;
L84 = 32'd631;
L85 = 32'd568;
L86 = 32'd618;
L87 = 32'd871;
L88 = 32'd827;
L89 = 32'd322;
L90 = 32'd1544;
L91 = 32'd1317;
L92 = -32'd413;
L93 = 32'd1214;
L94 = 32'd195;
L95 = -32'd610;
L96 = 32'd430;
L97 = 32'd1443;
L98 = 32'd193;
L99 = 32'd611;
L100 = 32'd476;
L101 = 32'd769;
L102 = 32'd1074;
L103 = 32'd1363;
L104 = 32'd1105;
L105 = 32'd435;
L106 = 32'd8;
L107 = 32'd492;
L108 = 32'd1587;
L109 = 32'd707;
L110 = 32'd1069;
L111 = -32'd209;
L112 = -32'd103;
L113 = 32'd69;
L114 = 32'd1428;
L115 = 32'd938;
L116 = 32'd236;
L117 = 32'd781;
L118 = -32'd20;
L119 = 32'd201;
L120 = 32'd122;
L121 = 32'd1050;
L122 = -32'd580;
L123 = 32'd1376;
L124 = 32'd2035;
L125 = 32'd1104;
L126 = 32'd959;
L127 = -32'd47;
L128 = -32'd32;
L129 = 32'd58;
L130 = 32'd425;
L131 = 32'd1460;
L132 = 32'd833;
L133 = 32'd291;
L134 = 32'd688;
L135 = -32'd431;
L136 = 32'd364;
L137 = 32'd446;
L138 = 32'd392;
L139 = 32'd1020;
L140 = 32'd486;
L141 = 32'd1185;
L142 = 32'd917;
L143 = 32'd16;
L144 = 32'd539;
L145 = 32'd872;
L146 = 32'd146;
L147 = 32'd483;
L148 = -32'd168;
L149 = 32'd175;
L150 = 32'd2200;
L151 = 32'd786;
L152 = 32'd1559;
L153 = 32'd2010;
L154 = 32'd254;
L155 = 32'd1160;
L156 = -32'd420;
L157 = 32'd781;
L158 = 32'd843;
L159 = 32'd822;
L160 = -32'd569;
L161 = 32'd413;
L162 = 32'd374;
L163 = -32'd0;
L164 = -32'd149;
L165 = 32'd991;
L166 = 32'd433;
L167 = 32'd523;
L168 = 32'd669;
L169 = 32'd92;
L170 = -32'd73;
L171 = 32'd53;
L172 = 32'd1254;
L173 = 32'd487;
L174 = 32'd1013;
L175 = 32'd715;
L176 = 32'd175;
L177 = 32'd731;
L178 = 32'd120;
L179 = -32'd263;
L180 = 32'd544;
L181 = 32'd502;
L182 = 32'd166;
L183 = 32'd664;
L184 = 32'd490;
L185 = 32'd741;
L186 = 32'd284;
L187 = 32'd831;
L188 = 32'd239;
L189 = 32'd908;
L190 = 32'd194;
L191 = 32'd1158;
L192 = -32'd11;
L193 = 32'd2031;
L194 = 32'd416;
L195 = 32'd315;
L196 = 32'd1578;
L197 = 32'd87;
L198 = 32'd1809;
L199 = 32'd1287;
L200 = 32'd1091;
L201 = 32'd882;
L202 = 32'd754;
L203 = -32'd124;
L204 = 32'd960;
L205 = 32'd552;
L206 = 32'd2231;
L207 = 32'd1000;
L208 = 32'd902;
L209 = 32'd661;
L210 = 32'd309;
L211 = 32'd1706;
L212 = 32'd152;
L213 = 32'd64;
L214 = 32'd1016;
L215 = -32'd212;
L216 = 32'd515;
L217 = 32'd175;
L218 = 32'd896;
L219 = 32'd878;
L220 = 32'd59;
L221 = 32'd716;
L222 = 32'd600;
L223 = 32'd410;
L224 = 32'd666;
L225 = 32'd44;
L226 = 32'd1306;
L227 = 32'd1349;
L228 = 32'd1451;
L229 = -32'd561;
L230 = 32'd1939;
L231 = -32'd211;
L232 = 32'd23;
L233 = 32'd1073;
L234 = 32'd158;
L235 = 32'd1435;
L236 = 32'd1131;
L237 = 32'd1059;
L238 = 32'd85;
L239 = 32'd1018;
L240 = 32'd621;
L241 = 32'd279;
L242 = -32'd153;
L243 = -32'd402;
L244 = 32'd385;
L245 = 32'd396;
L246 = 32'd672;
L247 = 32'd647;
L248 = 32'd451;
L249 = 32'd442;
L250 = 32'd590;
L251 = 32'd1141;
L252 = 32'd618;
L253 = 32'd734;
L254 = 32'd673;
L255 = 32'd302;
L256 = 32'd886;
L257 = 32'd612;
L258 = 32'd1107;
L259 = 32'd494;
L260 = -32'd178;
L261 = 32'd576;
L262 = 32'd1098;
L263 = 32'd1076;
L264 = 32'd1197;
L265 = 32'd2068;
L266 = 32'd507;
L267 = 32'd875;
L268 = 32'd935;
L269 = -32'd250;
L270 = 32'd680;
L271 = 32'd735;
L272 = 32'd1642;
L273 = 32'd1024;
L274 = 32'd899;
L275 = 32'd110;
L276 = 32'd566;
L277 = -32'd262;
L278 = 32'd771;
L279 = 32'd904;
L280 = 32'd81;
L281 = 32'd243;
L282 = 32'd1731;
L283 = 32'd361;
L284 = 32'd802;
L285 = 32'd183;
L286 = 32'd481;
L287 = 32'd1345;
L288 = 32'd358;
L289 = 32'd554;
L290 = 32'd1180;
L291 = -32'd913;
L292 = 32'd1027;
L293 = 32'd1224;
L294 = 32'd1461;
L295 = 32'd12;
L296 = 32'd1200;
L297 = -32'd71;
L298 = 32'd801;
L299 = 32'd1395;
L300 = 32'd1322;
L301 = 32'd1101;
L302 = 32'd895;
L303 = 32'd277;
L304 = 32'd868;
L305 = 32'd615;
L306 = 32'd468;
L307 = 32'd333;
L308 = 32'd924;
L309 = 32'd576;
L310 = -32'd276;
L311 = 32'd828;
L312 = -32'd604;
L313 = 32'd1286;
L314 = 32'd1077;
L315 = 32'd1879;
L316 = 32'd215;
L317 = 32'd4;
L318 = 32'd798;
L319 = 32'd923;
L320 = 32'd701;
L321 = 32'd707;
L322 = -32'd198;
L323 = 32'd913;
L324 = 32'd1479;
L325 = 32'd2275;
L326 = -32'd141;
L327 = 32'd1262;
L328 = 32'd565;
L329 = -32'd339;
L330 = 32'd679;
L331 = 32'd172;
L332 = 32'd308;
L333 = 32'd636;
L334 = 32'd1658;
L335 = 32'd1043;
L336 = 32'd643;
L337 = 32'd1486;
L338 = -32'd125;
L339 = -32'd410;
L340 = 32'd142;
L341 = 32'd396;
L342 = 32'd364;
L343 = 32'd377;
L344 = 32'd1225;
L345 = 32'd692;
L346 = -32'd471;
L347 = 32'd440;
L348 = 32'd761;
L349 = -32'd266;
L350 = 32'd1170;
L351 = 32'd205;
L352 = -32'd626;
L353 = 32'd1807;
L354 = 32'd446;
L355 = 32'd592;
L356 = -32'd51;
L357 = 32'd1393;
L358 = 32'd517;
L359 = 32'd78;
L360 = 32'd666;
L361 = 32'd1243;
L362 = -32'd82;
L363 = 32'd134;
L364 = 32'd604;
L365 = 32'd721;
L366 = 32'd560;
L367 = 32'd148;
L368 = 32'd214;
L369 = 32'd1456;
L370 = 32'd701;
L371 = 32'd1047;
L372 = 32'd984;
L373 = 32'd1010;
L374 = -32'd40;
L375 = 32'd803;
L376 = 32'd740;
L377 = 32'd1437;
L378 = 32'd366;
L379 = -32'd1012;
L380 = -32'd222;
L381 = 32'd158;
L382 = 32'd405;
L383 = -32'd568;
L384 = -32'd78;
L385 = 32'd320;
L386 = 32'd1575;
L387 = -32'd179;
L388 = 32'd1222;
L389 = 32'd232;
L390 = 32'd772;
L391 = 32'd835;
L392 = 32'd1114;
L393 = 32'd910;
L394 = 32'd928;
L395 = 32'd784;
L396 = 32'd1195;
L397 = 32'd1133;
L398 = 32'd936;
L399 = 32'd1049;
L400 = 32'd1377;
L401 = 32'd744;
L402 = 32'd63;
L403 = 32'd381;
L404 = 32'd932;
L405 = 32'd579;
L406 = 32'd993;
L407 = 32'd1046;
L408 = 32'd34;
L409 = 32'd814;
L410 = 32'd782;
L411 = -32'd60;
L412 = 32'd692;
L413 = 32'd1486;
L414 = -32'd476;
L415 = 32'd1061;
L416 = 32'd759;
L417 = 32'd385;
L418 = 32'd934;
L419 = -32'd250;
L420 = 32'd1061;
L421 = 32'd41;
L422 = 32'd522;
L423 = -32'd129;
L424 = 32'd118;
L425 = 32'd265;
L426 = 32'd1834;
L427 = -32'd19;
L428 = 32'd1330;
L429 = 32'd936;
L430 = 32'd763;
L431 = 32'd879;
L432 = 32'd1363;
L433 = -32'd117;
L434 = 32'd1368;
L435 = 32'd715;
L436 = 32'd157;
L437 = -32'd23;
L438 = 32'd803;
L439 = 32'd137;
L440 = 32'd388;
L441 = 32'd909;
L442 = 32'd752;
L443 = 32'd1084;
L444 = 32'd11;
L445 = 32'd829;
L446 = -32'd340;
L447 = -32'd674;
L448 = 32'd1521;
L449 = 32'd975;
L450 = 32'd225;
L451 = 32'd855;
L452 = -32'd400;
L453 = 32'd1732;
L454 = 32'd1100;
L455 = 32'd197;
L456 = 32'd1991;
L457 = -32'd358;
L458 = -32'd495;
L459 = 32'd687;
L460 = 32'd798;
L461 = 32'd244;
L462 = -32'd89;
L463 = 32'd163;
L464 = 32'd253;
L465 = 32'd670;
L466 = -32'd45;
L467 = 32'd532;
L468 = -32'd354;
L469 = 32'd1127;
L470 = 32'd433;
L471 = 32'd545;
L472 = 32'd124;
L473 = 32'd13;
L474 = 32'd603;
L475 = 32'd563;
L476 = -32'd202;
L477 = 32'd83;
L478 = 32'd451;
L479 = 32'd61;
L480 = 32'd1434;
L481 = 32'd410;
L482 = 32'd665;
L483 = 32'd589;
L484 = 32'd683;
L485 = 32'd785;
L486 = 32'd854;
L487 = 32'd636;
L488 = -32'd411;
L489 = 32'd722;
L490 = 32'd473;
L491 = 32'd160;
L492 = -32'd147;
L493 = 32'd742;
L494 = 32'd397;
L495 = 32'd156;
L496 = 32'd416;
L497 = 32'd577;
L498 = 32'd1525;
L499 = -32'd662;
L500 = 32'd842;
L501 = 32'd576;
L502 = 32'd851;
L503 = 32'd954;
L504 = 32'd338;
L505 = 32'd487;
L506 = 32'd1401;
L507 = -32'd107;
L508 = 32'd937;
L509 = -32'd141;
L510 = 32'd945;
L511 = -32'd26;
L512 = 32'd822;
L513 = 32'd795;
L514 = 32'd1481;
L515 = 32'd787;
L516 = 32'd992;
L517 = 32'd87;
L518 = -32'd54;
L519 = 32'd589;
L520 = 32'd49;
L521 = 32'd297;
L522 = 32'd1045;
L523 = 32'd240;
L524 = 32'd1244;
L525 = 32'd985;
L526 = 32'd1539;
L527 = 32'd356;
L528 = 32'd1128;
L529 = 32'd631;
L530 = -32'd178;
L531 = -32'd268;
L532 = 32'd1702;
L533 = 32'd1350;
L534 = 32'd706;
L535 = 32'd1371;
L536 = 32'd1439;
L537 = 32'd1522;
L538 = 32'd83;
L539 = 32'd746;
L540 = 32'd968;
L541 = 32'd1984;
L542 = 32'd1087;
L543 = 32'd791;
L544 = 32'd770;
L545 = 32'd221;
L546 = 32'd616;
L547 = 32'd1235;
L548 = 32'd450;
L549 = 32'd1035;
L550 = 32'd41;
L551 = 32'd1216;
L552 = 32'd1082;
L553 = 32'd1025;
L554 = 32'd109;
L555 = 32'd301;
L556 = 32'd1205;
L557 = 32'd1794;
L558 = 32'd5;
L559 = -32'd50;
L560 = 32'd644;
L561 = 32'd1221;
L562 = 32'd405;
L563 = 32'd832;
L564 = -32'd596;
L565 = 32'd292;
L566 = 32'd441;
L567 = 32'd451;
L568 = 32'd1408;
L569 = 32'd1604;
L570 = -32'd282;
L571 = 32'd1;
L572 = 32'd649;
L573 = 32'd975;
L574 = 32'd2247;
L575 = 32'd1671;
L576 = 32'd1089;

#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
#5
$display("%h", P);
$display("%h", P);

$finish;
end
endmodule
